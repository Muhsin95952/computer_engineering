module carry(C, A, B);
input A, B;
output C; 

and a1(C, A, B);
endmodule
