module not_gate(I, O);
input I;
output O;

not n_gate(O, I);

endmodule
