module buffer(I, O);
input I;
output O;

buf b_gate(O, I);

endmodule

