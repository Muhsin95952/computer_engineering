module andgate(I1,I2,O);
input I1;
input I2;
output O;

and a_gate(O,I1, I2);
endmodule

