module sum(S, A, B);
input A, B;
output S;

xor x1(S, A, B);

endmodule
