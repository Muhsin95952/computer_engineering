module MUX4x1_tb()
reg [3:0]I;
reg [1:0]sel;
wire out

MUX4x1 mymux(I, sel, out)

initial begin


