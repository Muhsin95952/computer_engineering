module MUX8x1_using_4x1_tb();
reg S0, S1, S2;
reg [7:0]I;
wire Out;

MUX8x1_using_4x1 c0(Out, S0, S1, S2, I);

initial begin
S0 = 0; S1 = 0; S2 = 0;
I[0] = 1; I[1] = 0; I[2] = 0; I[3] = 0; I[4] = 0; I[5] = 0; I[6] = 0; I[7] = 0;
#10
S0 = 0; S1 = 0; S2 = 1;
I[0] = 0; I[1] = 1; I[2] = 0; I[3] = 0; I[4] = 0; I[5] = 0; I[6] = 0; I[7] = 0;
#10
S0 = 0; S1 = 1; S2 = 0;
I[0] = 0; I[1] = 0; I[2] = 1; I[3] = 0; I[4] = 0; I[5] = 0; I[6] = 0; I[7] = 0;
#10
S0 = 0; S1 = 1; S2 = 1;
I[0] = 0; I[1] = 0; I[2] = 0; I[3] = 1; I[4] = 0; I[5] = 0; I[6] = 0; I[7] = 0;
#10
S0 = 1; S1 = 0; S2 = 0;
I[0] = 0; I[1] = 0; I[2] = 0; I[3] = 0; I[4] = 1; I[5] = 0; I[6] = 0; I[7] = 0;
#10
S0 = 1; S1 = 0; S2 = 1;
I[0] = 0; I[1] = 0; I[2] = 0; I[3] = 0; I[4] = 0; I[5] = 1; I[6] = 0; I[7] = 0;
#10
S0 = 1; S1 = 1; S2 = 0;
I[0] = 0; I[1] = 0; I[2] = 0; I[3] = 0; I[4] = 0; I[5] = 0; I[6] = 1; I[7] = 0;
#10
S0 = 1; S1 = 1; S2 = 1;
I[0] = 0; I[1] = 0; I[2] = 0; I[3] = 0; I[4] = 0; I[5] = 0; I[6] = 0; I[7] = 1;

end

initial
$monitor("S0 = %b S1 = %b S2 = %b I0 = %b I1 = %b I2 = %b I3 = %b I4 = %b I5 = %b I6 = %b I7 = %b Out = %b",
 S0, S1, S2, I[0], I[1], I[2], I[3], I[4], I[5], I[6], I[7], Out);

endmodule



